module Five_vote(A,B,C,D,E,Y);
	input A,B,C,D,E;
	output Y;
	reg Y;
	always @(A,B,C,D,E,Y)
		case({A,B,C,D,E})
		5'b00000:Y<=1'b0;
		5'b00001:Y<=1'b0;
		5'b00010:Y<=1'b0;
		5'b00011:Y<=1'b0;
		5'b00100:Y<=1'b0;
		5'b00101:Y<=1'b0;
		5'b00110:Y<=1'b0;
		5'b00111:Y<=1'b1;
		5'b01000:Y<=1'b0;
		5'b01001:Y<=1'b0;
		5'b01010:Y<=1'b0;
		5'b01011:Y<=1'b1;
		5'b01100:Y<=1'b0;
		5'b01101:Y<=1'b1;
		5'b01110:Y<=1'b1;
		5'b01111:Y<=1'b1;
		5'b10000:Y<=1'b0;
		5'b10001:Y<=1'b0;
		5'b10010:Y<=1'b0;
		5'b10011:Y<=1'b1;
		5'b10100:Y<=1'b0;
		5'b10101:Y<=1'b1;
		5'b10110:Y<=1'b1;
		5'b10111:Y<=1'b1;
		5'b11000:Y<=1'b0;
		5'b11001:Y<=1'b1;
		5'b11010:Y<=1'b1;
		5'b11011:Y<=1'b1;
		5'b11100:Y<=1'b1;
		5'b11101:Y<=1'b1;
		5'b11110:Y<=1'b1;
		5'b11111:Y<=1'b1;
		default:Y<=1'b0;
		endcase
endmodule