module CDEC(CS,LEDR1,LEDR2,LEDL1,LEDL2,SCOREAC,SCOREBC,RESULT);
	input [2:0]CS;
	output LEDR1,LEDR2,LEDL1,LEDL2;
	output SCOREAC,SCOREBC,RESULT;
	reg LEDR1,LEDR2,LEDL1,LEDL2;
	reg SCOREAC,SCOREBC,RESULT;
	always @(CS)
		case (CS)
			3'B000  :begin LEDR1<=1'B0;LEDR2<=1'B0;LEDL1<=1'B0;LEDL2<=1'B0;
						    SCOREAC<=1'B0;SCOREBC<=1'B0;RESULT<=1'B0; end
			3'B001  :begin LEDR1<=1'B1;LEDR2<=1'B0;LEDL1<=1'B0;LEDL2<=1'B0;
							SCOREAC<=1'B0;SCOREBC<=1'B0;RESULT<=1'B0; end
			3'B010  :begin LEDR1<=1'B0;LEDR2<=1'B0;LEDL1<=1'B1;LEDL2<=1'B0;
							SCOREAC<=1'B0;SCOREBC<=1'B0;RESULT<=1'B0; end
			3'B011  :begin LEDR1<=1'B0;LEDR2<=1'B0;LEDL1<=1'B0;LEDL2<=1'B0;
							SCOREAC<=1'B1;SCOREBC<=1'B0;RESULT<=1'B0; end
			3'B100  :begin LEDR1<=1'B0;LEDR2<=1'B0;LEDL1<=1'B0;LEDL2<=1'B0;
							SCOREAC<=1'B0;SCOREBC<=1'B1;RESULT<=1'B0; end
			3'B101  :begin LEDR1<=1'B0;LEDR2<=1'B0;LEDL1<=1'B0;LEDL2<=1'B0;
							SCOREAC<=1'B0;SCOREBC<=1'B0;RESULT<=1'B1; end
			3'B110  :begin LEDR1<=1'B0;LEDR2<=1'B1;LEDL1<=1'B0;LEDL2<=1'B0;
							SCOREAC<=1'B0;SCOREBC<=1'B0;RESULT<=1'B0; end
			3'B111  :begin LEDR1<=1'B0;LEDR2<=1'B0;LEDL1<=1'B0;LEDL2<=1'B1;
							SCOREAC<=1'B0;SCOREBC<=1'B0;RESULT<=1'B0; end
			default :begin LEDR1<=1'B0;LEDR2<=1'B0;LEDL1<=1'B0;LEDL2<=1'B0;
							SCOREAC<=1'B0;SCOREBC<=1'B0;RESULT<=1'B0; end
		endcase
endmodule 