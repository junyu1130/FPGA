module DCD7SG(A,LED);
	input [3:0]A;
	output [6:0]LED;
	reg [6:0]LED;
	always @(A)
		case(A)
			4'B0000 :LED <=7'B0111111;
			4'B0001 :LED <=7'B0000110;
			4'B0010 :LED <=7'B1011011;
			4'B0011 :LED <=7'B1001111;
			4'B0100 :LED <=7'B1100110;
			4'B0101 :LED <=7'B1101101;
			4'B0110 :LED <=7'B1111101;
			4'B0111 :LED <=7'B0000111;
			4'B1000 :LED <=7'B1111111;
			4'B1001 :LED <=7'B1101111;
			4'B1010 :LED <=7'B1110111;
			4'B1011 :LED <=7'B1111100;
			4'B1100 :LED <=7'B0111001;
			4'B1101 :LED <=7'B1011110;
			4'B1110 :LED <=7'B1111001;
			4'B1111 :LED <=7'B1110001;
			default :LED <=7'B1110001;
		endcase
endmodule